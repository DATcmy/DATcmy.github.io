��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  ��9�    LED�G���ެO����V��      �  ��_�    �@��1.5V���q������GLED      �  9QG    ���LED����      �  � 9G    ����LED����<      �  q 9� G    ����LED����<      �  9 ��    `�ߧ@���G�]�p�@�q���A�ϥΥ|�Ӷ}���H����l�����k�����A�Ϩ��l�@�e�Ჾ�ʤΥ��k��ʡA�q���u�i�Τ@��      �  	 a)o    l�ߧ@�T�G�ݧ�Ф����T�����ܿO�ΥH�ХܤT�Ӥ��P���A�@�@���T�a�Υs���ݧ�A�@�]�p�@�q���Ϭݧ��T�����ӳ��I��      �  1 y� �    �H��ݧ�i�����T�a      �  �i�w    <�ߧ@�|�G�ϥΤ@�ӹq���A��Ӷ}���A�]�p�@�q���������ʪ���V      �  �	 S     V�ߧ@�G�G�@���v��줺���U�@���A�ΩШⶡ�A�@�]�p�@�q�������k�A�@�ϦU�B���O�w�i�U�۶}��      �  9 	 )     c�ߧ@�@: �]�p�@�q���ϸ����εo���G����(LED)�@����w���U�ɵo�X�n���εo���A�@�����}���w���n���Υ��G����          �  �    ���  CLED_G�� 	 CTerminal  @TAi     :        "@���s�+�@  �  PTQi     <           ���s�+��    9$YT       
 ����    ��  CLED_Y�  � L� a     A        "@4֬q�@  �  � L� a     D           4֬q��    � � L       
 ����    ��  CLED�  0 L1 a     C        "@Ĳ��R��@  �  @ LA a     E           Ĳ��R���    ) I L       
 ����    �� 
 CBattery9V��  CDummyValue  h�h�    9V            "@      �? V �  h�i�      <           ���s�+�@  �  @�A�      :        "@���s�+��    ,�~      %    ��   �  !�#�  � �� �    9V            "@      �? V �  � �� �      D           4֬q�@  �  � �� �      A        "@4֬q��    � ��       )    ��   �  !�#�  X �X �    9V            "@      �? V �  X �Y �      E           Ĳ��R��@  �  0 �1 �      C        "@Ĳ��R���     �n       -    ��   �  !�#�  P�P�    9V            "@      �? V �  P�Q�      F          �r��{��=  �  (�)�      G        "@r��{���    �f`     1    ��   �  !�#�  ����    9V            "@      �? V �  ����      I    ���y�=?Ĳ��R��@  �  ����      H  �O�; "@Ĳ��R���    ���`     5    ��   �  ��  ����     H  �O�; "@Ĳ��R��@  �  ����     I    ���y�=?Ĳ��R���    �\��     8  
 ����    ��  0�1�     F          �r��{���  �  @�A�     G        "@r��{��=    )\I�     ;    ����    ��  @lA�     >         @8���ד@  �  PlQ�     ?        �8���ד�    9<Yl     >  
 ����    ��   l�     ;          �L�a㧝Խ  �  l�     @         �?L�a㧝�=    �<l     A    ����    ��  �l��     B         �?t�C��W>  �  �l��     9          �t�C��W�    �<�l     D    ����    ��  CBattery#�  p�p�    1.5V            �?      �? V �  p4qI     =         �?����ד�  �  p�q�      ?        �8���ד@    `��4    I    ��   �  F�#�  @�@�    1.5V            �?      �? V �  @�A�      >         @8���ד�  �  @4AI     =         �?����ד@    0�P4     M    ��   �  F�#�   � �    1.5V            �?      �? V �   4I     @         �?L�a㧝Խ  �   ��      ;          �L�a㧝�=    ��4    Q    ��   �  F�#�  ����    1.5V            �?      �? V �  ����      B         �?t�C��W�  �  �4�I     9          �t�C��W>    ���4     U    ��   �  ��  CSPDT��  CToggle  *�<      X  �  8d9y     `          �          �  XdYy     c          �          �  xdyy     d                       *:�d     [    ����P    ��  CMotorEM�  ����      7          �          �  �$�9     0          �          �� 	 CMechTerm       �                    \             �	�    3 	        �            ��$     `    ��  D `  bK�6�>       ���?<k<               ���?<k<W�Y�  � 4      d  �  �\�q     b          �          �  �\�q     _                     �  �\�q     ^          �            �2 \     f    ����P    W�Y�  � � 4      i  �  � \� q     5          �          �  � \� q     2          �          �  � \� q     ]                       � 2� \     k    ����P    ^��   �!�      \          �          �   �!     4          �          b�       �                    \             d�i�    8 	        �            �d�     o   ��  D `  bK�6�>       ��3X�#A               ��3X�#AW�Y�  �  D     r  �  � l� �     Y          �          �  � l� �     a                     �  � l� �     6          �            � Bl     t   ����P    !�#�  P �P �    9V            "@      �? V �  P �Q �      Z          �          �  ( �) �      [        "@             �f 0     y    ��   �  ��  CBuzzer�  �0�E      U          �          �  ����     X          �            �D�     }    ��  6 `  ��  ��1     S          �          �  ��1     W          �            ���     �    ����    ��  ()1     Q          �          �  891     *          �            !�A     �    ����    ��  CSPSTY�  � 0T     �  �  � |� �     O                     �  � |� �     /          �            � R|     �   ����P    !�#�  x �x �    9V            "@      �? V �  x �y �      .          �          �  P �Q �      N        "@            < �� �     �    ��   �  ��Y�  � �0�      �  �  � �� �     P          �          �   ��     -          �            � �0�     �    ����P    ��Y�  R���      �  �  `�a�     R          �          �  ����     ,          �            R���     �    ����P    ��Y�  ��8�      �  �  ����     +          �          �  �	�     )          �            ��8�     �    ����P    ��  1     V          �          �  ()1     T          �            �1     �    ����    !�#�  ����    9V            "@      �? V �  ����      o                     �  ����              "@            ����     �    ��   �  W�Y�  2���      �  �  @�A�     n          �          �  `�a�               �          �  ����                            2���     �    ����P    W�Y�  
�h�      �  �  ��     r          �          �  8�9�               �          �  X�Y�     p                       
�h�     �    ����P    ^��  ��      q   �~i8�*T`���Xw*  �  �|��     s   ��Ngm�K�T`���Xw�  b���PC.            1å*    \             ��     	 ��PC.    1å*    ��|     �   ��  D `  bK�6�>��PC.�DOGA�����а)��PC.�DOGA��Y�  �8 P\       �  �   � �      f          �          �   � !�      g          �            �Z P�      �    ����P    ��Y�  z8 �\       �  �  �� ��      i          �          �  �� ��                �            zZ ��      �    ����P    ��Y�  8 `\       �  �  � �                �          �  0� 1�                �            Z `�      �    ����P    !�#�  �� ��     9V            "@      �? V �  �� ��                 �          �  �� ��       e        "@            |� �@     �    ��   �  �� 	 CFilament#�          1W            �?      �? W �  �                �          �  d y     h          �            � d     �      ��`   ��#�  � �     1W            �?      �? W �  � �!     j          �          �  � !     k          �            �� �8     �      ��`   ��#�   �  �     1W            �?      �? W �  � %�      l          �          �  �� ��      m          �            $� �     �      ��`   ��  Xd Yy      L          �          �  hd iy                �            Q4 qd      �    ����    �� 	 CPushMake��  CKey  ( "@       �  �  l 	�      J          �          �  l �                �            � > !l      �    ����    !�#�  � � � �     9V            "@      �? V �  � � � �                            �  � � � �               "@            � � � @     �    ��   �  {��  �� ��       M          �          �  ��!     K          �            |� �     �    ��  6 `      �  �    ���  CWire  hhi�      < ݀  Phii     < ݀  @hA�      : ݀  � `� �      D ݀  � `� a     D ݀  � `� �      A ݀  @ �Y �     E ݀  @ `A �      E ݀  0 `1 �      C ݀  ����      H ݀  ����     I ݀  ����      I ݀  (�)�      G ݀  �)�     G ݀  P�      G ݀  PQQ     G ݀  PPQ�      G ݀  @�Q�     G ݀  0�1�      F ݀  0�Q�     F ݀  P�Q�      F ݀  pHqi      = ݀  @hqi     = ݀  @HAi      = ݀  p�q�      ? ݀  P�q�     ? ݀  @�A�      > ݀   Hi      @ ݀   hi     @ ݀  �i      @ ݀  ��     @ ݀   ��      ; ݀  �H�i      9 ݀  �h�i     9 ݀  ���i      9 ݀  ����     9 ݀  ����      B     �  �    �    �  �        �  �      �   �   �   �   �     � % � % & � & ) � ) * � * - � - . � . 1 � 1 2 � 2 5 � 5 6 � 6 8 8 � 9 9 � ; ; � < < � > > � ? ? � A A � B B � D D E E I I � J � J M � M N N � Q Q � R � R U U V V � [ [   \ \   ] ]   `   ` a a   c c   f f   g g   h h   k k   l l   m m   o   o p p   q q   t t   u u   v v   y   y z   z }   } ~ ~   � �   � �   � �   � �   � �   � �   �   � �   � � �   � �   � �   � �   � �   � �   � �   � �   �   � �   � � �   � �   � �   � �   � �   � �   �   � � �   � �   � �   � �   � �   � �   � �   � �   �   � �   � �   � � �   �   � � �   �   � � �   � �   � �   � �   � �   �   � �   � �   � � �   � %  �  & � )  �  * � -   �  . 8 6 9 � � 5 � 2 � � � � � � � � < � ; � � � � 1 I � � � N � � J ? � > M Q � � � � � B � A R V � �  � E  D U  t �        �$s�        @     +        @            @    "V  (      �                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 